module rettangolo(
//Posizione del rettangolo dall'angolo alto a sinistra
input [10:0] X_POS,
input [10:0] Y_POS,
//Controllo
input [10:0] X_CONTROLLO,
input [10:0] Y_CONTROLLO,

output CONFERMA
);

parameter altezza = 50;
parameter larghezza = 50;

//if (X_CONTROLLO > X_POS)

endmodule
